module dut_wrapper();
	initial
	begin
		$display("**DUT WRAPPER**BEGIN**");
		$display("**DUT WRAPPER**END**");
	end
endmodule
